library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity state_machine is
		port(
			X,Y, CLK: in std_logic; -- Inputs
			Z: Out std_logic
		);
end state_machine;

Architecture behave of state_machine is
------------------- 00. STATE DEFINITIONS -------------------
	signal state: integer range 0 to 3:= 0;



begin	-- beggining the behavioral portion or architecture
------------------- 01. STATE REGISTER -------------------
	process(CLK) -- setting up the clock
		begin
			if(CLK'event and CLK='1') then
				case state is
				-- directions for the 0 state
				when 0 => if X='0' and Y='0' then state <= 0;
  		        elsif X='0' and Y='1' then state <= 1;
				elsif X='1' and Y='0' then state <= 2;
				elsif X='1' and Y='1' then state <= 1;
				end if;

				-- directions for the 1st state
				when 1 => if X='0' and Y='0' then state <= 1;
        		elsif X='0' and Y='1' then state <= 0;
				elsif X='1' and Y='0' then state <= 2;
				elsif X='1' and Y='1' then state <= 3;
 				end if;

				-- directions for the 2nd state
				when 2 => if X='0' and Y='0' then state <= 2; 
        		elsif X='0' and Y='1' then state <= 3;
				elsif X='1' and Y='0' then state <= 3;
				elsif X='1' and Y='1' then state <= 1;
				end if;

				-- directions for the 3rd state
				when 3 => if X='0' and Y='0' then state <= 3; 
        		elsif X='0' and Y='1' then state <= 0;
				elsif X='1' and Y='0' then state <= 1;
				elsif X='1' and Y='1' then state <= 0;
				end if;
			
			end case;
		end if;
	end process;



------------------- 03. OUTPUT LOGIC -------------------
Z <= '1' when (state = 2) or (state = 3) else '0';

end behave;
